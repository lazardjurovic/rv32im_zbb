class bram_sequencer extends uvm_sequencer#(bram_seq_item);

endclass : bram_sequencer