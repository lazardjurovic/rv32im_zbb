`ifndef AXI_SEQ_PKG_SV
`define AXI_SEQ_PKG_SV

    import uvm_pkg::*;      // import the UVM library
    `include "uvm_macros.svh" // Include the UVM macros

    `include "axi_seq_item.sv"
    `include "axi_sequencer.sv"
    `include "axi_base_seq.sv"
    `include "axi_transaction.sv"
    `include "axi_read_stop_flag.sv"
    `include "axi_reset_low_seq.sv"
 
`endif
