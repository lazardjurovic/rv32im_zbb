`ifndef CONFIGURATION_PKG_SV
 `define CONFIGURATION_PKG_SV

   import uvm_pkg::*;      // import the UVM library   
 `include "uvm_macros.svh" // Include the UVM macros

`include "cpu_config.sv"


`endif
