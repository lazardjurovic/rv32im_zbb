class cpu_scoreboard extends uvm_scoreboard

endclass : cpu_scoreboard